`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   18:20:03 10/07/2016
// Design Name:   rrefs
// Module Name:   C:/Users/User/Desktop/Processor-20161003T064542Z/rrefs/tb.v
// Project Name:  rrefs
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: rrefs
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb;

	// Inputs
	wire [31:0]inv11;
	wire [31:0]inv12;
	wire  [31:0]inv13;
	wire  [31:0]inv14;
	wire [31:0]inv15;
	wire  [31:0]inv21;
	wire  [31:0]inv22;
	wire  [31:0]inv23;
	wire  [31:0]inv24;
	wire  [31:0]inv25;
	wire  [31:0]inv31;
	wire  [31:0]inv32;
	wire  [31:0]inv33;
	wire  [31:0]inv34;
	wire  [31:0]inv35;
	wire  [31:0]inv41;
	wire  [31:0]inv42;
	wire  [31:0]inv43;
	wire  [31:0]inv44;
	wire  [31:0]inv45;
	wire  [31:0]inv51;
	wire  [31:0]inv52;
	wire  [31:0]inv53;
	wire  [31:0]inv54;
	wire  [31:0]inv55;

	// Instantiate the Unit Under Test (UUT)
	rrefs uut (
		.inv11(inv11), 
		.inv12(inv12), 
		.inv13(inv13), 
		.inv14(inv14), 
		.inv15(inv15), 
		.inv21(inv21), 
		.inv22(inv22), 
		.inv23(inv23), 
		.inv24(inv24), 
		.inv25(inv25), 
		.inv31(inv31), 
		.inv32(inv32), 
		.inv33(inv33), 
		.inv34(inv34), 
		.inv35(inv35), 
		.inv41(inv41), 
		.inv42(inv42), 
		.inv43(inv43), 
		.inv44(inv44), 
		.inv45(inv45), 
		.inv51(inv51), 
		.inv52(inv52), 
		.inv53(inv53), 
		.inv54(inv54), 
		.inv55(inv55)
	);

	initial begin
		// Initialize Inputs
		

	end
      
endmodule

